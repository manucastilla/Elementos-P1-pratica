------------------------------
-- Elementos de Sistemas
-- Avaliacao Pratica 1
--
-- 10/2019
--
-- Questão 2 - Seven Seg
------------------------------

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity sevenSeg is
  port (
    H : in  STD_LOGIC_VECTOR(3 downto 0);
    a,b,c,d,e,f,g : out STD_LOGIC );
end entity;

architecture  rtl OF sevenSeg IS


begin



end architecture;
