corsi@corsi-note.26690:1568381085